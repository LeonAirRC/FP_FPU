library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity sub_inner is
    port (
        num_a : in std_logic_vector(31 downto 0);
        num_b : in std_logic_vector(31 downto 0);
        output: out std_logic_vector(31 downto 0);
    );
end sub_inner;

architecture arch_sub_inner of sub_inner is



begin



end architecture;